module abc (in1,in2,out);
input in1,in2;
output out;
and a1 (out,in1,in2);
//assign out = in1 & in2;
endmodule